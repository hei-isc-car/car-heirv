ARCHITECTURE studentVersion OF hb_gen IS
BEGIN

  hb <= '1';

END ARCHITECTURE studentVersion;
